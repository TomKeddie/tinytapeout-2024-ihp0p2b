`default_nettype none

module uart_tx (
                input  clk,
                input  reset,
                output tx_pin0,
                output tx_pin1,
                output tx_pin2,
                output tx_pin3,
                output tx_pin4,
		output tx_pin5
                );

  wire [7:0]           text0 [0:49];
  wire [7:0]           text1 [0:49];
  wire [7:0]           text2 [0:49];
  wire [7:0]           text3 [0:49];
  wire [7:0]           text4 [0:49];
  wire [127:0]	       text5 [0:68];
   

  // a couple of random things to push out a serial port
  assign text0[0]  = "T";
  assign text0[1]  = "i";
  assign text0[2]  = "n";
  assign text0[3]  = "y";
  assign text0[4]  = "T";
  assign text0[5]  = "a";
  assign text0[6]  = "p";
  assign text0[7]  = "e";
  assign text0[8]  = "o";
  assign text0[9]  = "u";
  assign text0[10] = "t";
  assign text0[11] = " ";
  assign text0[12] = "I";
  assign text0[13] = "H";
  assign text0[14] = "P"; 
  assign text0[15] = " ";
  assign text0[16] = "0";
  assign text0[17] = "p";
  assign text0[18] = "2";
  assign text0[19] = " ";
  assign text0[20] = "N";
  assign text0[21] = "o";
  assign text0[22] = "v";
  assign text0[23] = "2";
  assign text0[24] = "0";
  assign text0[25] = "2";
  assign text0[26] = "4";
  assign text0[27] = " ";
  assign text0[28] = "T";
  assign text0[29] = "o";
  assign text0[30] = "m";
  assign text0[31] = "K";
  assign text0[32] = "e";
  assign text0[33] = "d";
  assign text0[34] = "d";
  assign text0[35] = "i";
  assign text0[36] = "e";
  assign text0[37] = " ";
  assign text0[38] = " ";
  assign text0[39] = " ";
  assign text0[40] = " ";
  assign text0[41] = " ";
  assign text0[42] = " ";
  assign text0[43] = " ";
  assign text0[44] = " ";
  assign text0[45] = " ";
  assign text0[46] = " ";
  assign text0[47] = " ";
  assign text0[48] = "\r";
  assign text0[49] = "\n";
  
  assign text1[0] = "O";
  assign text1[1] = "p";
  assign text1[2] = "e";
  assign text1[3] = "n";
  assign text1[4] = " ";
  assign text1[5] = "t";
  assign text1[6] = "h";
  assign text1[7] = "e";
  assign text1[8] = " ";
  assign text1[9] = "p";
  assign text1[10] = "o";
  assign text1[11] = "d";
  assign text1[12] = " ";
  assign text1[13] = "b";
  assign text1[14] = "a";
  assign text1[15] = "y";
  assign text1[16] = " ";
  assign text1[17] = "d";
  assign text1[18] = "o";
  assign text1[19] = "o";
  assign text1[20] = "r";
  assign text1[21] = "s";
  assign text1[22] = ",";
  assign text1[23] = " ";
  assign text1[24] = "H";
  assign text1[25] = "A";
  assign text1[26] = "L";
  assign text1[27] = " ";
  assign text1[28] = " ";
  assign text1[29] = " ";
  assign text1[30] = " ";
  assign text1[31] = " ";
  assign text1[32] = " ";
  assign text1[33] = " ";
  assign text1[34] = " ";
  assign text1[35] = " ";
  assign text1[36] = " ";
  assign text1[37] = " ";
  assign text1[38] = " ";
  assign text1[39] = " ";
  assign text1[40] = " ";
  assign text1[41] = " ";
  assign text1[42] = " ";
  assign text1[43] = " ";
  assign text1[44] = " ";
  assign text1[45] = " ";
  assign text1[46] = " ";
  assign text1[47] = " ";
  assign text1[48] = "\r";
  assign text1[49] = "\n";

  assign text2[0]  = "I";
  assign text2[1]  = "'";
  assign text2[2]  = "m";
  assign text2[3]  = " ";
  assign text2[4]  = "s";
  assign text2[5]  = "o";
  assign text2[6]  = "r";
  assign text2[7]  = "r";
  assign text2[8]  = "y";
  assign text2[9]  = ",";
  assign text2[10] = " ";
  assign text2[11] = "D";
  assign text2[12] = "a";
  assign text2[13] = "v";
  assign text2[14] = "e";
  assign text2[15] = ".";
  assign text2[16] = " ";
  assign text2[17] = "I";
  assign text2[18] = "'";
  assign text2[19] = "m";
  assign text2[20] = " ";
  assign text2[21] = "a";
  assign text2[22] = "f";
  assign text2[23] = "r";
  assign text2[24] = "a";
  assign text2[25] = "i";   
  assign text2[26] = "d";
  assign text2[27] = " ";
  assign text2[28] = "I";
  assign text2[29] = " ";
  assign text2[30] = "c";
  assign text2[31] = "a";
  assign text2[32] = "n";
  assign text2[33] = "'";
  assign text2[34] = "t";
  assign text2[35] = " ";
  assign text2[36] = "d";
  assign text2[37] = "o";
  assign text2[38] = " ";
  assign text2[39] = "t";
  assign text2[40] = "h";
  assign text2[41] = "a";
  assign text2[42] = "t";
  assign text2[43] = ".";
  assign text2[44] = " ";
  assign text2[45] = " ";
  assign text2[46] = " ";
  assign text2[47] = " ";
  assign text2[48] = "\r";
  assign text2[49] = "\n";

  assign text3[0]  = "Y";
  assign text3[1]  = "o";
  assign text3[2]  = "u";
  assign text3[3]  = " ";
  assign text3[4]  = "a";
  assign text3[5]  = "r";
  assign text3[6]  = "e";
  assign text3[7]  = " ";
  assign text3[8]  = "i";
  assign text3[9]  = "n";
  assign text3[10] = " ";
  assign text3[11] = "a";
  assign text3[12] = " ";
  assign text3[13] = "m";
  assign text3[14] = "a";
  assign text3[15] = "z";
  assign text3[16] = "e";
  assign text3[17] = " ";
  assign text3[18] = "o";
  assign text3[19] = "f";
  assign text3[20] = " ";
  assign text3[21] = "t";
  assign text3[22] = "w";
  assign text3[23] = "i";
  assign text3[24] = "s";
  assign text3[25] = "t";
  assign text3[26] = "y";
  assign text3[27] = " ";
  assign text3[28] = "p";
  assign text3[29] = "a";
  assign text3[30] = "s";
  assign text3[31] = "s";
  assign text3[32] = "a";
  assign text3[33] = "g";
  assign text3[34] = "e";
  assign text3[35] = "s";
  assign text3[36] = ",";
  assign text3[37] = " ";
  assign text3[38] = "a";
  assign text3[39] = "l";
  assign text3[40] = "l";
  assign text3[41] = " ";
  assign text3[42] = "a";
  assign text3[43] = "l";
  assign text3[44] = "i";
  assign text3[45] = "k";
  assign text3[46] = "e";
  assign text3[47] = ".";
  assign text3[48] = "\r";
  assign text3[49] = "\n";

  assign text4[0]  = "T";
  assign text4[1]  = "e";
  assign text4[2]  = "d";
  assign text4[3]  = " ";
  assign text4[4]  = "P";
  assign text4[5]  = "a";
  assign text4[6]  = "r";
  assign text4[7]  = "k";
  assign text4[8]  = "e";
  assign text4[9]  = "r";
  assign text4[10] = " ";
  assign text4[11] = "2";
  assign text4[12] = "3";
  assign text4[13] = " ";
  assign text4[14] = "M";
  assign text4[15] = "a";
  assign text4[16] = "r";
  assign text4[17] = " ";
  assign text4[18] = "1";
  assign text4[19] = "9";
  assign text4[20] = "4";
  assign text4[21] = "2";
  assign text4[22] = " ";
  assign text4[23] = "-";
  assign text4[24] = " ";
  assign text4[25] = "1";
  assign text4[26] = "2";
  assign text4[27] = " ";
  assign text4[28] = "A";
  assign text4[29] = "p";
  assign text4[30] = "r";
  assign text4[31] = " ";
  assign text4[32] = "1";
  assign text4[33] = "9";
  assign text4[34] = "9";
  assign text4[35] = "5";
  assign text4[36] = " ";
  assign text4[37] = " ";
  assign text4[38] = " ";
  assign text4[39] = " ";
  assign text4[40] = " ";
  assign text4[41] = " ";
  assign text4[42] = " ";
  assign text4[43] = " ";
  assign text4[44] = " ";
  assign text4[45] = " ";
  assign text4[46] = " ";
  assign text4[47] = " ";
  assign text4[48] = "\r";
  assign text4[49] = "\n";

assign text5[ 0 ] = 128'b00000000000001111111111111110110001111110001111111001111111111111111111001111011000111101001011111111111111111100111000000000000;
assign text5[ 1 ] = 128'b00000000110100111111111111111101100011111100011111100011111111111111111110111111110011111010000111111111111111110111111100000000;
assign text5[ 2 ] = 128'b00000000111101000111111111111110011000111111000111111001111111111111111010000111111100111101110001111111111111111101111111000000;
assign text5[ 3 ] = 128'b00000110001111010011111111111111100110001111110001111111111111111111111111110001111110001111011100111111111111111111011111110000;
assign text5[ 4 ] = 128'b00001101100111110100111111111111111011000011111100011111111111111111111111111011010111100011110100101111111111101111111111111000;
assign text5[ 5 ] = 128'b00011011010001111010001111111111111110110001111111001111111100111111111111111110100111111000111101111011111111111011111111111100;
assign text5[ 6 ] = 128'b01010010111100011110100011111111111111101100011111110011111111011111111111110111100011111110001111010101111111111110111111111110;
assign text5[ 7 ] = 128'b10011111111011000111101000111111111111111011000111111000111111010111111101111111010000111111100110110111111111111111111111111111;
assign text5[ 8 ] = 128'b10101110001110110001111010001111111111111100110001111110000000000000000000001001010100001111110001101011111110101111111011111001;
assign text5[ 9 ] = 128'b11101011100111111100011110100011111111111111001100000000000000000000000000000000000100100011111100011011111111101111111100111110;
assign text5[10 ] = 128'b11111110110101111111001111101001111111111111100000000000000000000000000000000000000000011101111111000110101111111010111111011111;
assign text5[11 ] = 128'b11111100111100011111100011110110011111111100000000000000000000000000000000000000000000000100101111110001111111111111101111110110;
assign text5[12 ] = 128'b11111111111011000111111000111101000111100000000000000011111111111111111111111000000000000000011111111100010111111111110011111101;
assign text5[13 ] = 128'b11101111110100110001111110001111011110000000000000111111101011010001111111111111110000000000000101101111001101101101110100111111;
assign text5[14 ] = 128'b01111011111101001000011111100011111000000000000111111001111110101100011010111111111110000000000001010111100011010111011101011111;
assign text5[15 ] = 128'b01111100111111010110001111111011100000000000111111111111111011101011000110101011111111110000000000011101111000110101110111010111;
assign text5[16 ] = 128'b11001111011111100101100011111110000000000011111111111111101110001010110001011010011111111100000000001111011110001111011111110101;
assign text5[17 ] = 128'b11110011110111111001011000111100000000001000111111001111111011100101101100110100111111111111100000000011011111100011110111111111;
assign text5[18 ] = 128'b01111100111101111110110111111000000000000000000000000000000000000000000000001101101111111111110000000001011111111000111101001111;
assign text5[19 ] = 128'b10111111001111011111101111100000000000000000000000000000000000000000000000100011010111101111111100000000111111111110011111011101;
assign text5[20 ] = 128'b00101111100011100111111111000000000000000000000000000000000000000000000000001000110110111111111110000000001101111111100111111110;
assign text5[21 ] = 128'b10011111111010111001111110000000000000000000000000000000000000000000000000011110001101111111111111000000001011111111110001111111;
assign text5[22 ] = 128'b11000111111110011110111100000000000000000000000000000000000000000000000000110101100010110111111111110000000101101111111100011111;
assign text5[23 ] = 128'b11110001111111100111111100000000000000000000000000000000000000000000000000011111011001101101111111111000000010111011111111000111;
assign text5[24 ] = 128'b11111100011111111111111000000000000000000000000000000000000000000000000000110110110110011011111111111000000001100110101111110001;
assign text5[25 ] = 128'b00111111000110111111111111111111111111111111111100000000000001111111111001011101101111000110101111111100000000001000111111111100;
assign text5[26 ] = 128'b01110111110011111111111111111111111111111111111100000000000001111111111110100101011010110001101011111110000000110011000001111110;
assign text5[27 ] = 128'b10010101101100111111100000000111111111011111111100000000000000110111111111101101100110101100011011111110000000111101101110011111;
assign text5[28 ] = 128'b10101001011010001111000000001101111111110111111100000000000001101110111111111010011011101011000101111111000000011111011111101111;
assign text5[29 ] = 128'b11001001010100101111100000001111011111111111111100000000000000111011101111111101101111111110110001111111000000011111110111111001;
assign text5[30 ] = 128'b11110011100101111111100000001011111111111111111100000000000000000000000000000000000000000000001000111111000000011111111101111000;
assign text5[31 ] = 128'b11111101111011011111000000011110111101111111111100000000000000000000000000000000000000000000000010011111000000011111111111111110;
assign text5[32 ] = 128'b11111111011111111111000000000111101110011111111100000000000000000000000000000000000000000000000001111111100000001101111111111111;
assign text5[33 ] = 128'b01111110010101111111100000011101110011100111111100000000000000000000000000000000000000000000000101011111000000000111111111111111;
assign text5[34 ] = 128'b11011111101111011111100000011110110001111011111100000000000000000000000000000000000000000000000011011111000000010111111111111111;
assign text5[35 ] = 128'b11110111111011111111100000000111101001011111111100000000000000000000000000000000000000000000000001111101000000011100111111111111;
assign text5[36 ] = 128'b11111001111110111111100000000001111111110111111100000000000000000000000000000000000000000000000011111111000000011111001111111111;
assign text5[37 ] = 128'b11111110011111111111100000001100011111100111111100000000000001111111100000000000001111111111111111111110000000011111110011111111;
assign text5[38 ] = 128'b11100111101111111111110000000011001111111011111100000000000001111111100000000000001111111111111111111111100000000111111100111111;
assign text5[39 ] = 128'b10101001111011111111110000000110110011111011111100000000000000111111100000000000000011111111111111111100000000110001111111011111;
assign text5[40 ] = 128'b11101110111100111111111000000001001000111111111100000000000001111111100000000000000100111111111111111100000000101100011111100111;
assign text5[41 ] = 128'b01111011111011101111111000000001011010001111111100000000000001011111100000000000001011011111111111111000000011011011001111111001;
assign text5[42 ] = 128'b00011110110111110111111100000000110101100011111111111111111111111111100000000000001010100011111111110000000001110111100011111100;
assign text5[43 ] = 128'b11001111101101011111111110000000000101011000101101111011111111111111100000000000000110101001111111100000000110101111111000111111;
assign text5[44 ] = 128'b10100011011111000111111111000000001011111110011011011000111111111111100000000000000001101011111111000000001111111111111110001111;
assign text5[45 ] = 128'b11111000110101110101111111100000000011110011100110110110111111111111100000000000001100010110111100000000011111111110011111100011;
assign text5[46 ] = 128'b11110110001101011111111111110000000001111001010001111011101111111111100000000000001111001101111000000000111111111111000111111000;
assign text5[47 ] = 128'b01011101100011010111111111111000000000011011101100011110011111111111100000000000000111100011100000000011111111111111110011111110;
assign text5[48 ] = 128'b10011111011000101101111111111110000000000100101011000111101110011111100000000000000101111110000000000111111111111111111100111111;
assign text5[49 ] = 128'b11100111110110011011011111111111000000000001010010110001111011111111100000000000000001011000000000010111111111111111111110001111;
assign text5[50 ] = 128'b11111001111001000110101100111111110000000000000011111100111110111111100000000000000011100000000001110100111111111111111111100011;
assign text5[51 ] = 128'b11111110111111010001101111111111111100000000000001111111001111111111100000000000001111100000000000111111001111111111111111111000;
assign text5[52 ] = 128'b11111111101111101100011000111111111111100000000000000111110011111111100000000000001111000000011110011111110011111111111111111110;
assign text5[53 ] = 128'b11111111111111111011000111101101111111111000000000000000000000111111100000000000001111000001111111000111111100011111111111111111;
assign text5[54 ] = 128'b11111111111110101110110001111010011111111111000000000000000000000000000000000000001111001110001111110001111110000111111111111111;
assign text5[55 ] = 128'b11111111111111101111101100111110111111111111111100000000000000000000000000000000001111101111100111111100011111100011111111111111;
assign text5[56 ] = 128'b11111111111111110111011010001111111111111111111111111000000000000000000000000001111111111011110000111111000111111000111111111111;
assign text5[57 ] = 128'b11111111111111111101110110100011110111111110111111111111111111111110011111110010111111111111111100011111110001111110001111111111;
assign text5[58 ] = 128'b00111111111111111111111101011000111101110011111111111111111111101111100111101000111111111111001111000111111100111111100011111111;
assign text5[59 ] = 128'b10001111111111111111110111010110001111011010111101111110111110001011110001111010110111111111110011110001111110001111111000111111;
assign text5[60 ] = 128'b00100011111111111111111111110111100011110110101111011111101111100010111100011110100001111111111101111100011111100011111100011111;
assign text5[61 ] = 128'b01011000111111111111111111111011111001111101110111101111111011111000101111000111101010011111111111011111000111111000111111111010;
assign text5[62 ] = 128'b00110100001111111111111111001110111100011011111000111100111100111110010111110011111010010111111111110111100111111110001111111100;
assign text5[63 ] = 128'b00011101001111111111111111110111101111000110111100011100001111001111100101111100111110000001111111111101111110111001100011111000;
assign text5[64 ] = 128'b00001111010001111111111111111100001011110001101111010111011111110111110111011110001111010000111111111110011111001011111001110000;
assign text5[65 ] = 128'b00000011110101011111111111111111000010111100011011111101111111111101111100010111100011110100001111111111100111101110111100000000;
assign text5[66 ] = 128'b00000000111101011111111111111011111111101111000101111111011111111111111111010101111000111101001011111111111011100011101100000000;
assign text5[67 ] = 128'b00000000000110100111111111111100111101110111110011011111000111111111110111110001011110001111011101111101111110111101000000000000;

   wire [7:0]	       char_space = " ";
   wire [7:0] char_at = "@";
  reg [3:0]            bit_counter;
  reg [5:0]            text_index;
  
  reg                  tx_pin0_int;
  reg                  tx_pin1_int;
  reg                  tx_pin2_int;
  reg                  tx_pin3_int;
  reg                  tx_pin4_int;
  reg                  tx_pin5_int;
  assign tx_pin0 = tx_pin0_int;
  assign tx_pin1 = tx_pin1_int;
  assign tx_pin2 = tx_pin2_int;
  assign tx_pin3 = tx_pin3_int;
  assign tx_pin4 = tx_pin4_int;
  assign tx_pin5 = tx_pin5_int;

  always @(posedge clk) begin
    // if reset, set counter to 0
    if (reset) begin
      bit_counter <= 0;
      tx_pin0_int  <= 1'b1;
      tx_pin1_int  <= 1'b1;
      tx_pin2_int  <= 1'b1;
      tx_pin3_int  <= 1'b1;
      tx_pin4_int  <= 1'b1;
      tx_pin5_int  <= 1'b1;
      text_index   <= 6'b0;
    end else begin
      // bit counter - START, 8xDATA, STOP, IDLE = 11 bits
      if (bit_counter == 10) begin
        // reset
        bit_counter    <= 0;
         if (text_index == 49) begin
          text_index <= 6'b0;
        end else begin
          text_index <= text_index + 1;
        end
      end else begin
        // increment counter
        bit_counter <= bit_counter + 1;
      end
      case(bit_counter)
        0       : begin
          tx_pin0_int = 1'b1; // idle
          tx_pin1_int = 1'b1; // idle
          tx_pin2_int = 1'b1; // idle
          tx_pin3_int = 1'b1; // idle
          tx_pin4_int = 1'b1; // idle
          tx_pin5_int = 1'b1; // idle
        end
        1       : begin
          tx_pin0_int = 1'b0; // start
          tx_pin1_int = 1'b0; // start
          tx_pin2_int = 1'b0; // start
          tx_pin3_int = 1'b0; // start
          tx_pin4_int = 1'b0; // start
          tx_pin5_int = 1'b0; // start
        end
	9       : begin
          tx_pin0_int = 1'b0; // upper bit
          tx_pin1_int = 1'b0; // upper bit
          tx_pin2_int = 1'b0; // upper bit
          tx_pin3_int = 1'b0; // upper bit
          tx_pin4_int = 1'b0; // upper bit
          tx_pin5_int = 1'b0; // upper bit
	end
        10      : begin
          tx_pin0_int = 1'b1; // stop
          tx_pin1_int = 1'b1; // stop
          tx_pin2_int = 1'b1; // stop
          tx_pin3_int = 1'b1; // stop
          tx_pin4_int = 1'b1; // stop
          tx_pin5_int = 1'b1; // stop
        end
        default : begin
          tx_pin0_int = text0[text_index][bit_counter-2];
          tx_pin1_int = text1[text_index][bit_counter-2];
          tx_pin2_int = text2[text_index][bit_counter-2];
          tx_pin3_int = text3[text_index][bit_counter-2];
          tx_pin4_int = text4[text_index][bit_counter-2];
          tx_pin5_int = char_at[bit_counter-2];
        end
      endcase
    end
  end
endmodule
